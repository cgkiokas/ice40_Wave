FunctionGen_pll_inst: FunctionGen_pll
port map(
          REFERENCECLK => ,
          PLLOUTCOREA => ,
          PLLOUTCOREB => ,
          PLLOUTGLOBALA => ,
          PLLOUTGLOBALB => ,
          RESET => 
        );
